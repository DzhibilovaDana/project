module GreenP (
	
	// pins for FPGA
	inout M1,
	inout P3,
	inout T7,
	inout T6,
	inout T5,
	inout T4,
	inout T3,
	inout T2,
	inout P2,
	inout N2,
	inout L2,
	inout K2,
	inout J2,
	inout G1,
	inout F1,
	inout C2,
	inout D3,
	inout E5,
	
	inout N5,
	inout N3,
	inout R7,
	inout R6,
	inout R5,
	inout R4,
	inout R3,
	inout R1,
	inout P1,
	inout N1,
	inout L1,
	inout K1,
	inout J1,
	inout G2,
	inout F2,
	inout B1,
	inout D4,
	inout D5,

	//pins for periphery
	inout T14,
	inout R13,
	inout T13,
	inout R11,
	inout M10,
	inout P9,
	inout N9,
	inout M9,
	inout M8,
	inout N8,
	inout P8,
	inout N12,
	inout M11,
	inout T11,
	inout R10,
	inout T10,
	inout R9,
	inout T9,
	inout T8,
	inout R8,
	inout N6,
	
	inout C16,
	inout B12,
	inout A12,
	inout B11,
	inout A11,
	inout B9,
	inout A9,
	inout A8,
	inout B8,
	inout A7,
	inout B7,
	inout A6,
	inout B6,
	inout C6

);

    assign N9 = G1;

    assign M9 = N5;
endmodule